library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package CHESS_TYPES is
    type boardType is array(63 downto 0) of integer range -6 to 6;
    type colorMatrixRev is array(399 downto 0) of natural range 0 to 3;
    type colorMatrix is array(0 to 399) of natural range 0 to 3;
    
constant letterG : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,0,
0,0,0,1,1,1,1,1,1,1,1,1,1,1,2,0,0,0,0,0,
0,0,3,1,1,1,1,1,1,1,1,1,1,1,1,2,0,0,0,0,
0,0,3,1,1,3,3,3,3,3,3,3,1,1,1,1,2,0,0,0,
0,0,3,1,1,2,0,0,0,0,0,0,3,1,1,1,1,2,0,0,
0,0,3,1,1,2,2,2,2,0,0,0,0,3,1,1,1,2,0,0,
0,0,3,1,1,1,1,1,1,2,0,0,0,3,1,1,1,2,0,0,
0,0,3,1,1,1,1,1,1,2,0,0,0,3,1,1,1,2,0,0,
0,0,0,3,1,1,1,1,2,0,0,0,0,3,1,1,1,2,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,3,1,1,1,2,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,3,1,1,1,2,0,0,
0,0,0,2,2,0,0,0,0,0,0,0,0,3,1,1,1,2,0,0,
0,0,3,1,1,2,0,0,0,0,0,0,0,3,1,1,1,2,0,0,
0,0,3,1,1,1,2,2,2,2,2,2,2,1,1,1,1,2,0,0,
0,0,3,1,1,1,1,1,1,1,1,1,1,1,1,1,2,0,0,0,
0,0,0,3,1,1,1,1,1,1,1,1,1,1,1,2,0,0,0,0,
0,0,0,0,3,1,1,1,1,1,1,1,1,1,2,0,0,0,0,0,
0,0,0,0,0,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterA : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,3,3,3,3,3,3,0,0,0,0,0,0,0,
0,0,0,0,0,0,2,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,0,0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,2,2,2,2,1,1,1,3,0,0,0,0,
0,0,0,0,2,1,1,3,0,0,0,0,2,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,3,3,3,3,3,2,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,3,2,2,2,2,2,2,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterM : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,3,3,3,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,
0,2,1,1,1,3,0,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,2,1,1,1,1,3,0,0,0,0,0,0,2,1,1,1,1,3,0,
0,2,1,1,1,1,1,3,0,0,0,0,2,1,1,1,1,1,3,0,
0,2,1,1,1,1,1,1,3,0,0,2,1,1,1,1,1,1,3,0,
0,2,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,3,0,
0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,
0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,
0,2,1,1,1,3,1,1,1,1,1,1,1,1,2,1,1,1,3,0,
0,2,1,1,1,3,2,1,1,1,1,1,1,2,2,1,1,1,3,0,
0,2,1,1,1,3,0,2,1,1,1,1,2,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,2,1,1,2,0,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,0,2,2,0,0,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,2,1,1,1,3,0,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,0,2,2,2,0,0,0,0,0,0,0,0,0,0,2,2,2,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterE : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,3,3,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,2,2,2,2,2,2,2,2,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,3,3,3,3,3,3,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,2,2,2,2,2,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterO : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,2,2,2,2,2,2,1,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,1,3,3,3,3,3,3,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterV : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,3,3,3,3,0,0,0,0,0,0,0,0,3,3,3,3,0,0,
0,2,1,1,1,1,3,0,0,0,0,0,0,2,1,1,1,1,3,0,
0,2,1,1,1,1,3,0,0,0,0,0,0,2,1,1,1,1,3,0,
0,2,1,1,1,1,3,0,0,0,0,0,0,2,1,1,1,1,3,0,
0,2,1,1,1,1,1,3,0,0,0,0,2,1,1,1,1,1,3,0,
0,0,2,1,1,1,1,3,0,0,0,0,2,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,3,0,0,2,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,3,0,0,2,1,1,1,1,1,3,0,0,
0,0,0,2,1,1,1,1,3,0,0,2,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,3,2,1,1,1,1,1,3,0,0,0,
0,0,0,0,2,1,1,1,1,3,2,1,1,1,1,3,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,0,0,2,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,0,0,0,0,2,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,1,3,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterR : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,2,2,2,2,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,3,3,3,3,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,3,3,3,3,1,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,2,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,2,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,2,2,0,0,0,0,0,0,0,2,2,2,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterW : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,0,0,0,0,0,0,0,0,0,3,3,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,0,3,3,3,0,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,3,0,2,1,1,1,3,0,2,1,1,1,3,0,
0,0,2,1,1,1,1,3,1,1,1,1,1,3,1,1,1,1,3,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,0,0,2,1,1,1,1,1,2,1,1,1,1,1,3,0,0,0,
0,0,0,0,0,2,1,1,1,2,0,2,1,1,1,3,0,0,0,0,
0,0,0,0,0,0,2,2,2,0,0,0,2,2,2,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterH : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,0,0,0,0,0,0,0,0,3,3,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,3,3,3,3,3,3,3,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,3,2,2,2,2,2,2,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,0,2,2,2,0,0,0,0,0,0,0,0,2,2,2,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterI : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,0,2,2,2,1,1,1,3,3,3,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,2,2,2,1,1,1,3,3,3,0,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,0,2,2,2,2,2,2,2,2,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterT : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,2,2,2,2,1,1,1,3,3,3,3,3,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterB : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,3,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,2,2,2,2,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,3,3,3,3,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,3,2,2,2,2,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,3,3,3,3,3,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterL : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,2,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterC : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,0,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,2,2,2,2,2,2,1,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,2,2,2,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,0,3,3,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,0,3,1,1,1,3,0,0,
0,0,2,1,1,1,1,3,3,3,3,3,3,1,1,1,1,3,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,0,0,0,2,2,2,2,2,2,2,2,2,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterK : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,0,0,0,0,0,0,0,3,3,3,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,1,3,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,2,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,2,1,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,3,0,2,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,3,2,1,1,1,1,3,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,3,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,3,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,3,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,2,1,1,1,1,3,0,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,2,1,1,1,1,3,0,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,2,1,1,1,1,3,0,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,2,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,1,3,0,0,
0,0,0,2,2,2,0,0,0,0,0,0,0,2,2,2,2,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterN : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,3,3,3,0,0,0,0,0,0,0,3,3,3,0,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,3,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,3,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,3,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,3,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,3,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,2,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,2,1,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,2,1,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,2,1,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,2,1,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,2,1,1,1,3,0,0,0,0,0,2,1,1,1,3,0,0,0,
0,0,0,2,2,2,0,0,0,0,0,0,0,2,2,2,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant letterS : colorMatrix := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,3,0,0,0,0,
0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,2,2,2,2,2,2,2,2,2,2,0,0,0,
0,0,2,1,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,2,1,1,1,1,3,3,3,3,3,3,3,3,0,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,1,1,1,1,3,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,3,0,0,
0,0,0,3,3,3,3,3,3,3,3,3,3,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,
0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,
0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,
0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant pawnSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,1,2,2,2,2,2,2,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant rookSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,1,1,2,2,1,1,2,1,0,0,0,0,0,
0,0,0,0,0,1,1,0,0,1,1,0,0,1,1,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant knightSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,1,0,1,1,0,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,1,1,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,1,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,1,1,1,2,1,1,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant bishopSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant queenSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,1,1,2,2,1,1,2,1,0,0,0,0,0,
0,0,0,0,1,1,1,0,0,1,1,0,0,1,1,1,0,0,0,0,
0,0,0,0,1,0,0,0,0,1,1,0,0,0,0,1,0,0,0,0,
0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

constant kingSymbol : colorMatrixRev := (
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,1,2,2,2,2,2,2,2,2,2,2,1,0,0,0,0,
0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
0,0,0,0,0,0,1,2,2,2,2,2,2,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,1,2,2,2,2,1,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,1,1,1,2,2,1,1,1,0,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,1,2,2,2,2,2,2,2,2,1,0,0,0,0,0,
0,0,0,0,0,0,1,1,1,2,2,1,1,1,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,1,2,2,1,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
end package;